`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
PBxUhVrtWQEYOgb846Uv1sblkfb858tIOxXo5rSddtfNCCEaO6prOlrL6WWMok0v65NKAfNc24ct
xvcfwfVZn6pJLtI6aSJSRmTxG5GbjARcdFUpEQDBtUa4sAPMQtfZH1EIXufrcyxVW0XHTR7NfmbF
qvS0f84o1Ixfwgq0s4SVZ/cR5eixxcDOHJkeGNuRCF8c6r1aIEuE11tFlfos8wa2S7uhzhbhuAwd
jGnf13Ugn2l/BiuYbYpvg32KZvVGytJZ/jIKoOwtmjqDITZa9eS5uZFPmhCfqiaLfARe3gEdJwDM
VrP/j9Bw3m49r5kbYv/sPEvDIayVLCOr4ijwUA==
`pragma protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vG2MIsh9mK5WFqR7CZiQxAiJjbEpC8txbekQw6AfJ6/VWnF89geya0NQH3sioSl/yDNpWpXtEBqO
z8AJUbElhPqIDYzXPiEivSobyySonx2X0uCdcJouNl/v0FPaAQYCK8AUE3Ge2s3hse1XbmVqv7ZP
Y5qolN4zu0TOIlg4vB1+BTsuFow0v/IEoGR50X3yMj+DdCUIuRjl9OoX3lWT0rqw970MkQ5WOvn/
ZhsGOUVEa5swEGx5pTWK9rS4lS/s1q4YcLbS5OeSKnfTm7Bma4dQ3aKFmH4Jo37S3bHaAjADHSyc
OlA4EtFlsKlzzNfFcxoUhg7KfxitvBb2tophTw==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FV/3fpCT9rfkvj7vGf7H4iFLwONfv5yUkaBm4abp14Iadl/Ybdv2xjQOEAL0pWkfms08npBI7t4G
msUrfE93qg==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
iJhKydg23OP7sBpn7z4PB8q7WBOyQUXWMrIV2O/pWxlypf/RpKvTeWta7ZjeHIXrqYW1vATfnFYH
KffZziTGeXMp0GDONlIFq2Qla3fM1pmdSK3IvrPeNuYlsf+WfUT6uvjfunXWqXPT1fVLz7/0Nab1
ZnEsI4HXb/InsBjQim3VpKHPBlQeNERl9hExuvQYyS8r+j2mqTzgR+EES5zMdJJsUq6Tk6UGI5wF
d6kRUT5r5qEt50jaEfKFDj75HP1n7Tuasfr8O0MevqYvj98QmnFIDYepEkt9Ljvkvt/yj3gSID2M
4qrc/kttTD2TaB6JvKAqAO/Szpm3E9kRZBvB6A==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
TmA+sceFhlvNvYoL3GY2zygozlF2gKEQ4A5fIxzBaE0qXgC1YQhRjonQx+YYb5tG5J1TDYLtRBfS
v64j9USAdax/8kivVBMVXKqBBMqD+V2j1xsrLI8nng3HNOGBDyzpVrjQxPiBYmEwYm127I0k5tAB
q7f8Zcp5BA9A7YiPZVY=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
CtnoIChRHsmy/qBOvdecE+A1dR3wjyYuWKMfO1jOidf6ynMANArGWc4r8HTO7qhb1Z4TbmmEG89J
a0jZpsPvxqCpPRB0YoWCFbVuM3vxpRqy7OROD7ITd6q+0g8KOWanxPlLr6bT2HROZon50SO2azln
zb6EkIdjSMV8bP6d6M3SQlpW3rgtCkCmga5xhWGy0K8JOBPzJ7zD/GwwRrDPtnRR0DpyrDo1g8b2
l6QmdEomvQn6E8HRw0JKjEC23lGcNkXHWjFNLUO98cSrHh+H8o8nUdrw2qANJ9nJz6+xGN6t0T3f
m/EjUs3a4bAUqt01dDjnoiZuPVm0OJdsfBLJ0g==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
UrGwKDd/1QadwaGJuP8846x2A993ximCAJapb3bMaPSGBDEO9A0jPErFBA1KVOVeTK/6GREITCOO
kQUCBMGX84xmB3DKN/vtNJgs+hR53/RkssvaFt3utock0Fu3jmW6G8oAlZPUk5xuz3ZclLLk3zd7
b4+6GhssWTcJZUQTpFtfSHf9rzJtOVnfvssBzD9n9rKAavWOn0jgzU8w7LFG78jesOkkDRuf5AEC
O/3gMfhEbMgOvVlrw0VjgEMmnsmLjNJseq9mTu+TWFCtTTOhmTzkslcKwAqE5RGc85+QZ+Y7YTjh
vhXzh1hnBiJhadKuJFBNWiA0xJ7fT/yTmf0Jaw==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ZE+5HsZ7+s4D77YRJB7qciSuBMFSXam+Uezzo5KOHGOvuK0Czz+aZpjVDST9UUaxh5O+2DWaNkZd
K9zMBV9T+VTBgjlh7HzI5cbxtm+L7apsp+J2vwBKBmsNYO3LVgMnHYm+uECtR2dEfpGjFYUotmcX
ndknm7PwpJAlpEzkR0w=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
falKwGnr8t27uIOToebSrqeBQrBP5mPjpmoZpQ1b1QgLCIjb1Ax/qMTs0S0FkVIDlxDo0yuqRw1V
fyxzO19ZgTzsaVJCXVWZsRvnv3nCrJ7X74FSf7SUyvyEaBclCXZiqJSwHtK6tFrMBtfZiQQn+0of
l8weOHHNTljKfv+syccV4ZugkBMZ4Hj+YMWVAosOPpmJZZqhufSArsA3XzI4cR1HWHTSVcOPo6aj
c40rYyZrBcS9o/pXNBh4EgMfTFOYi2H7ye7r54YffFTwFKpy3qtNgZcOWFTiKY5yNG6DcPpT8hoP
xVSzIoXfxs+YszrfP7J1YsK4h3Evv0srY3RWtg==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
98pxjlvfQ9nOY2K4eowaSh8qTVmo7cno2cFtJKE60nCqSAm67p1pD2dsncHsWeGHjhbUvVmliH9y
TjFjBvqHUU0Fgev+82rjXG4k7LGAKNhrWWLr1qfSUQy6sUMlIPVcF8amdWWROGC7L10Txo7dN3HG
VONAfsV3hR1HPDyHj7/9u9rnAgiIRXf2sdmCBh65Lp9ATKMo0Yxtaq5vxw7aJbc7lkagLWzMLlDB
pWRWqI2Yi30QkAtQJI5ii0sKIjScjg0lBrnlgBR/T8A6DdO2KYZRvEUQMB5pmNvTjWvU+a87/qsd
r3/7/chpJIjsmvWiGHFhMc4tBjB8823K3Mt/N5xgMYvCsUHzN1IOpbaVM8K92bkY1vrYf+I6o52b
6MoFrsnwZKVyKv944Q8F14DRrog8TbD6D8lWG15DgJn/YZSZ98pDFY77OtYswNdp9YzSS+clJlHh
VJHz1NbO7p0TcDpm6+Pb4MpbMPaaVZ8zGsRi/BvP0UcVi2ORZDfL6snLZgfR1yLqNU++buaytkwE
tyR6SZO4aU6iAAprLsy5Lil9qDuR8h1z/M7T4B0Q2WDAcCgJ52fdnHoSwcUmXEcf3k6MD/xJTEHn
disnxyKEoJqcDrbU674ESWLz4/Y96p2riNm7R+wXNb1zDIWg2iiAJsTIUgleGM7+AEj5HcULSR2u
zxhmMcII5D8YnnxIkFrUwXXjAhUjsJ4edt25CBpIF1oG8iq2H72LBxLie0IPNV9WzAJyQR6gkaT8
QhAIz/n/e3WQFSqjJfIhXozTVlx5WeB3lawLk04ZjipyQ4JSH5vTS3Jwm/gBH5plYyLI6o7vIrIr
bhRFdsfYVJw+5i2+AkUtXq0c8ne8bQPqym24LuFVEmgy/0EwbHKUsSb0sKfrdOhJk5cj6GDX7Xhk
7qUhHFXpHnrN4A5h4BBrKOe8RWt0KzanYeR4xabnjgHrYvUo93cT1WwL5nO6kvJHy+n4nE1OHfyg
vuTN/jsfhgCva1wBb4XsPYcfGVorTUqGXw3RmAWSXmW/gHG4He1mRE3NvayAZvIyCn7XNAAaH5Q8
zLjIjjwjisohTcbehvH6dMZoPvGhB+9/p5WaaKNSqKTBoop1pqa2Y5QCCzDyS5R/BI2Cf7AbgmE6
i7GgVAYVytNdoIQrLdCmtKL89d4ORmZjF2ibyEWClAuw6BkZZFPHB2ZQZa7V0qY7g8l5xZc/KHni
zebKwjBnTx8Vmhm/DJm0GE8Wo3XIgce4+8SL1jKR8gq2zacLlKKune1xKAwyJNdGoFueJAUDhsTT
Q5T8uG+PUF7R8c6pmyLLQfnS7nYZGtflGrKazvxWYl7HF9kGGm61X2UwENZRTDAskq8xRf4TrJR3
xTLiEP5YpJTChPiDr9ZJ3YRsGj8sdrDYLJHVuyEN1pW+vLxKZTkzsbnfwj2cSwtGlBk+tKztc40H
2i4OKt6uuKKfvUEkIXwlM59uSTaGSXy56M7yT3lrokuEdZ/aX4jNarYwgMmlYifL4vtur2OYKNZ4
Fg4qQJO9HkXFzFpgf8TZr5OUpFAljCfdeV892U0ajcUisO/ZQ/bmgunycR07xGZRBeiSp7nw+rSG
6AxeXSRXGKtyCXrPhsibLV99pZR2c6an+HF0697qz3BZW0zahpHIYv9wV1iuQM7x2hMEuDUes3DL
MIYrxGSx+mBqeEiyNAmmTcm5btIGx8kqtLHL6zUYd8vhvqqXCNVxHhnXFGJLAZN4Mddrq5E/IvcS
ZU7M569VF+xlL7BlRbcY6XNJqtmDm6HBUGPukBHW2rQMtddVU0kpkSGZZiFzB354zea8nOqTy7fG
XzEfXm1eVUNaAamH11r1S1vFQPX9bBL86jAIaTTTBsMySqlLd+Oc35N2KAuQfSbqWx4tYQmJO2YK
8+gbiyr2q+tfsfOlsyKsKV8XgD52XKFAPQAWSB5PRNP+wJx0iR97gZdixp9ES/Uj6FGIDSr7LFY6
oURxIPPFPPt9SmdO2n8EsuDMHS0UqUL5YC2xgP9rQYQNxf/W/vwK8DyoWS3J7GiZtOcu6orXDF4g
zQ4ZOJhtfNPnMH7JU7URpEr2uAi0lZxitQ31UqwqH1z3Jfawl3HFXfDJi1I2mVfk/6HDdvADNImA
/rTmvkAdBHlIVYeq9UpSPMiAdoj+59Si2iDESwzhQbGMbpHj1qVo00AF3DgsEQtbA3EuR2fmnYgx
sG9VHg2awLNn5mPP+BBCRqUJ9M6DmQ9LttJ8cuJKVB/x5uOzwr/Q4DzsswTdfmIRUKjBecldxI90
dLZvZ4hv8hbKWfM+mdzPyNowFGFTP3XHxxXTiY1cLDmCbfCQaC4aJFXFHWTnI2avExHTcg9r4v1m
Xf9V72+bm9NoYjX01Gzn4NsmIZGA5yA0yabZJ0kEiE6xW/2WVYJWC+FV5ZjV/ChLGehQhoCxepO9
UogViDp3qwmHi/GEUXIJ82gK+peX73Fj8/MWBnNNwzsWXRo0/RQWR74Z3PryQrO4U5w90XYu8Xc/
+yFW2vs5BXh/4p8l+Ycchj2BKM9l5rwT+bOwYE7tVkcnOnBVnIuipeeUrNsUUltYTJuL8L2BF7fT
USjaZhmxWX+CBP9tiEjSnEq4b4EoNpU7VU3mt5e2NR548Kj1TQ43MpwbB7YAcsEro+frIBn05D93
eMysGV6rGAfLp33w+nq7X2Rk26oQ0Fj6HR3ADzK8IZPBBqCuJJEucNjjx4Syfj4YIznh6Z5+IIqh
fD6ZmJDbkybZocad8cIBrPYBONVAu7msYZRQFgng4GiVa617bdUwz1zVMSpWZ3q3j64baqXuWoVv
pcBfHuCzTGsAc+xLngFLNNih2DpChYIANkRbRQAuRGWqFlaHmA25O5fWyyXhkxDrbcRpg82Y2Udq
qE1lg70Fz/mJ+rkoQT1RNmj5WsDr4oJDph9ykR8tIpZH+bHS7xt4rUEo4m1PrJsHh6LmdDcwOGFS
7JcZWbPwqb/JjMafCMTZ4TCquHb8GINs5sxwCaJ/dh6EjdPvw2Dv69TkZsJlxXjHjybzeRLq8DMy
VYAkt0oO53Ri+FHNbHM1VgTLysXMcJe/woD0OPwmPwwg4a5GVa6NwWU/6SHHYF6VaHz402qI4edC
3LArYJ3UU3fesUcucnV5WAVXusxvEPOgVw0zOmrFlBaXnFBjkczQ1+aH7JB3FJEeITwwpJp8h2jE
MzwkLHerKQtjWHnShzBMD6K3+BgSRc+bdRZRBPBvJSeopMa5c7YT9vhD/vTe2IZp79MZYhiG1an9
AbRjrj/hrqAzC+iCOxDXGjefTY9CsCoO9Z0ERZG+xfebITdquLuO3qoYeYGT83mbsdUAdmkzcyTb
m3SqbUiJCZjeR0KaJ5o5Wl5iN/Jolx+lswfsVutoLAdLXnf96HYPgS2zSKQs6zuXHdbPAu3nCX/H
/Cn0RSExjt5VeL3240v28qsTqkXefLj2MpQs0qtblloyXViaw19qbwj1iQMAMYHrwA7zCpqi9XJW
pPSELBnA7MVUB20m+0TuiGYYfXVojrOe0LRd+tTW2pZKw6O/j0/1tiN8jG2EpJf/H1r2eoqRJ3O0
J1I9LlgU+kXJMyT/9NOloy7mDoOrP26Y/f5k35+OZc1lld9PRANgn4K36u6nukcKjtQf/HiUasoZ
rcRFAaCsRBpZixdFOArB9eBxPvwEXMz/WsDo0HY4quXR8os6ZLU0UAImhQa5jXqnYVP1vf6IPL/F
NerWWOG95iEI/Jgojq+sNusq8/KaC4vKRa2RBeXfUsHTwD5TaOrES5Cy6FwPl90fFmcX1oehijj0
hqzctn2yeNpkJSix/W0jTGCd4Pza+47E9xOo5osFrHKhJWVOMs91dikdONCgJ8Eb9KWzuTWW7Cz4
mgbWSa4z2x6eWXZCLJyC+etvElcctB4syKU9LXA3mRXtXJMze+X1zRZAPn+uXR8GLaqlzluKSkhV
os1rDxTC+s4hTkc8qGCBBt4B6SO0KQS8h505PIKRtbCAtvyvWoBCTK2RjEQdW4cn7VX4o8Cq6UOJ
OIQFdQWGs35vXpSGESRtZdXtY2NeLK3i4ix3wmMPf6qwHrYHfnkXEu0/OaGR+c7jX6Y1RubRlazB
oRSc9dMkvn2iA7hE4THjFWh5psWw0BEB65ul2vzPLUq4J8c54mVYbThe0hS5dBV6k11rZq5EmUUh
iYYatvs9HtIX6Q60RvcMbb3B+QprZbkqKSOOkmEx3B2WekL4gF++exwIXYoJK3dwvFsfWgaUWXOH
F3PV48HAuoSKBQS08Nue4bro9Pv8gpNWFZ5VEhJWDbtiv7YjMoC8UGoAMFPrNNN0lIfN4DYi5HRU
WXwqWnziwIyzj2G6JRygiHl7pw9TU9ZlVUR0pGjgm0qCwNljej3QMtSJPkZ+tjpu+DRYRqcZ1ADT
U3TVWXAxFuVyCqmblHqELuuCiE5emNWa/LPB38ho/0xs/6bLRYkBl6Q/qtKOt3jsEFYdoI0TFLuQ
j4FPac1nMLqdZSRjCUtZR1rer9tAmuEhUauUfI1sziRa6xQRAm6Atqx58ElSk0i4W6oQwRKpnOuk
sShbv8sQCK8vyUsmgbqLpW2lYCnAIE7wdyhr24QEegyYoW+cSLMZ+sU+tqatXZ/vgCPEtX0nzjZ9
WMGmixPWUP4dHyCLHjo8tWda59o3C4jtK/5GiBVH8ttuiuG6KWwfSPAw189HKoqZ3nRVKbnCukAu
MwCw5UaL5imxfjgebTt5Ecag+N2f0dTPgjACzrM9ZfrdbP1bKmWh5cT9NTn2A18Hk+NCnaMkiQ+j
nj3m/f++u/vgKTAqEp4NboRrL2SMT6eQ4muc84TLZ3ZKQ8j4WQAB6J0gZnvjgWr0UrmhKP9/RKcH
20v2zzDTQHE76SAGn/uamLq026Owb2deMxAvW8Q8eo0f2poD6S2pXmlr8co0osd2s6g5lVEzsb6U
JmOqpe1NvexpFdr8h0W1LIGWuZp0SjLe3oAI5ByBIvn+cG1unAmiS5qPszpQ6N84siZuhP+N/9HD
62y25DeQcR3qIJOnhALuO/YmpBAKp7WrHwyHvRYpp1bpYC1Fmbt65WoC+zE3PmKm0q3zBf4Tc6Vp
HCyxykhX52PIjdKhFKF6hOopb+CLyAjP9Il24QAIixXbPDPLA3aqZoNjP1k9/LLfS67agUCz4drM
S4oyUmo4lpx1mSKVuUeMgfUQBRAR2FmtBBkCKt19JcmyXPmKfQB5aeuKq1XqgNXtjCHsbgNSzAGN
kqRaftusoPW33JcgOJhWFB3DQ7WpaWIWcVJdomltrTa2osxqqzE/Uf1EbIiUMgoKKv+mj+IiKY7G
Bu/twY6TVhOY6KM171fTXh9JnmffaebMI3iHZlXC7ds71xg3pHE+ZTAAcXf/NopCnBnQoGueAkCe
63s75tRT2/ykCaC7TUnLMCd8iAxM5K29Xs7+wJz0WfR8cE5XQ/eR37GjHKRSxZQgpak8ahNEAMP0
A/NoJolnw+5Zgv5Yecc1sIWJS6J+zgwsGVw2bcKKpwRDlbM2VuSkRIEDhFgk50TXmtODHaLUTYlm
IiiPokfoSbzI7QQ34JOhMQ7U2EFpKw68L6E1CKhT8qvOuY6l2va1ccANPy8nUGzkYLs4yOLGQDfc
7DRQrXP7kPF4vJWKROHxRAlRDKaLT70tFliGcmo8IVnlYwLbbZJNdyLrrBww0gQQ5rLZVFH9mjEE
t0e7m6f1b4xEELUZij51ASP1NpG0aJgbkW85W1zuRSl0oFTeEeiUJguW3Cs0adN+FSGoutSmD9Ud
Bks9NN2uCp5C1TDpQFs4k2KqzST7NnRJy+9fytQpXW9LtcPlltROTAkmKH5ISacrYWYcGI/jMWcK
aRpt8uLAai3OuVHSG6QugmPj4y2KhVcpR3bzhp9Ka7QWMXLS3fC51/djm08Y3IaY0Wav91lh1Cho
1kDhSVCllSLgfv4W7+Mse7SKMewM918/g8cB1AQLIjfg2Fe/xdrM3uynP4G5RjsvXftXfH0tkGYO
rl0jtQzKjIQTkO+j8TvfKdcYJs+j9Dz1pYc8H0VSKsy9sEaVU5PEJcR0QNpeY4v/aPS2RZRJ4wip
iBlg3TLo5NMJKqtg9Wilfc2VlocG0YUXeoCGSS+p1WHC1PKqGE16V1PMId14hUlnAWHRZwEPfSmB
cyK+kXR/6vP2k5W7SmVLk5tmvcweCpTWArszdV0BgU58ZFFAMXI7MdZ4tXlEJ8iogdVDPpCJxI52
bS/xdWDAijQET/G0fkHDbhzUJZqJlSHeIYTVyr/f4EhMT2rUb9MwZhXJmLQ1p8EDjFrfvi4qAKTc
Bpe+hoH421nCImkvNbSmww6Tuha97C+flLbulKM/YjqupYRa5R/4k+T9oV37bpCfn28OZzf/IIPA
OAhzGdPTSH4yyrJLPR+nab7Ua1FzFhitYIfjaMQEBnmvCGk5b8K9JBHQOMMyhRbfzD3yFKBaI28/
OFOccWgIIao7/LCZ/qrk9thWPlmsROxkyfWdUzyIG6NQb05CXEM3vO82t8ZpVCuYXhpwvHWcX88K
V30LMePWEzDoKYN3Yfqd7TZUGi5dsgVW53q8R4NJByeWxYpnySAxkQlshtsEjGsq+n2xUw+C4jK0
AgaytaBVIaNoOXwLexGHWBKeXk2GkXTTCvKvSF9ZUNEPQL7tyjcmKdOe9V/VhVGBdp/yp0Wplhl2
1iO8TbXiwH0OO5/ttNKiaH2ouTzdv/u7Z52YBf/PTmlrd6z4j7RslXEDpOtkMpX1bl9dSyD4qgPC
EG4Y2Kj1GIRwg0g9lH1/It+wp+2rekmKKQy8jGzZDk5y6pdMHmv2erG58aQ39eVDjnPWiPYDfvL9
ZU+0CMeogA0T4Y45BEQyR6KJt6qJJ+A/vQ+xRSSk9a37q0oQ+ade7lLdnRojNkC/3hggk3FM54n8
TffXYAeYCip677V1++rBDbsoEANUcTKyKbEr4Z//g9Oiq3HG8xY6Jo6/OumWZQo9knpKnHnWc4ad
zuiGKLqg8PagNuI8p+4NjA7Kkq1TckfyWt4OFXGayTsXJwqvFwfVgth5kdDlCIP7gez9iwW0Zs/k
cFYNfCh2U8v71s6tQhzIs8t7LZgA+Vki3+3JixDsqfFdnLSSm/xFpJRu+TreTRNIisZrcFxzWdsR
V233ZGjoW2iUcM/DtiBJwZJeKCsDYGpk+0eELk/3uL5tkRv/n9zO9Noqd0jdH8sN0dTAF9PKU88T
d9W39DLTzpBHFBuFULux2xXPitABfkSPBYly+70tpVubvNx7kf7sPhPC7/Y0Z2pNRgGnR4UV2zGv
obtHcV71Jmk4X5YYZo6/8eElAkiGoSijIi5OjRH4yG8GIr+5jX5Tg/uAhvB+NoWZWgveUK+zgCJQ
pPLNooyxGPj6amrCDo+uPl+yTYQ1zBlHa7DIQb+GTC3i3URVNNiXbSY30TfUAWTpPjIBonfZ/z7N
Io3hE4xANoHDBk9s29yeKvr1oVsGl/mdv3YBAwzSa+Ti5t+8D+IttJyH4kN1fs03Hjhe8HgdhX+a
neaM+nsvS3+tALh64M516RbYS6wrlR4sdVUGOVczJyW3rR/tPrC9Si757Qypeb2iLN27T3e4tKBV
3zHsN+oifJfstaIsMs/dihgE3S8xRmU6zzjMlaP+rDzz3N0uF5aGqzchL8dUcJgtpjK6XwjPW8Ur
1v1YJE3226XQ1DVTP/0BN4srOk8mrT2en38SgILpLUAEEcIsChRcQ5JDhzmK4QtMcl0nKxHKKGWj
X3jPVQxfemDN3cuhUzldxY1o9LkuRjO1IXqrLsn0LmFc9AEoDVsurMvKUakFSYGHea1VhHVrYXW9
EsGz/BbirF/m8rdQDecpMLW6yM/IilSSm2yPljUhjH10AZyy5/ROeRt71Fi021DJT1dTTlU6WHBv
IWWIcUdvVq68BlwYM5QVdfsp7sB2Pfan1fDFWpoDLlNrFUjjKt/DfIog/0rpIGncddsV8K52AMcw
ofpJ+l7pCu6/aWetH4HWPaYvTyIDe04uQfEIdPOXJmA8o7Z0HiPGrUs57TvBzynd/LSGgISly6gt
9J9WFw/kD3EIDhIP8o8HuJ4/vUVC5isAlhl0d3APtoXULZvaE7x66JukU6oT2KFubLx15Q0emeV2
1+Vb5xpaDsfGd5Z9EZ2T5k0qC2jmu0IB+yuh0IVR8J7VJMGqWeaYHKyLCPk8xoKdEOWjte8NPc3D
0Ci9DLHaqZzdVShSzOZS7ga3lNqHDPG88Gm4r8+7eb2Hv4qbkJbZzLWuh8SsrjGzpGIzkXf5n8dH
eZ1vt8orDsObk7UT1o+w5Md6TRdPbanziJZ9+/W3KYZHsDZoxBYPS65ycnsUU+pL3bDNleBT277H
KLsO/kpLz3DvujD5N1iXJHYByhMtdiiS4dMCLWU9Vxce9otQGlKAULREZeaH5oIsOEn+POVH9m2+
a5BRiOA7NSPfOdN7+wLkb5lwq2sHaH8jRjycNwo9RwBFas/iwRnHaOCn+4jVke2QdAWCpKGc3eao
/SiABINOEsp2JJgTQp10Joefr+D/ZIcKdVQ+KlDi1bDIL9yzyVPQHZK81LegVERIWcjMROQ/Vdye
zgR3qxPt5ckJWIWBl3aLDDGZGvroLyDsn9ZzeAWgTLaBnxVAVm5UegHsSx1Nf/zM95Dmr+ny161k
eROdtrIZVKYNiLA9kBTo98OHlUaDpixAfcLvSGRHEAsieiJCNeROIIHK5BxfcGUrCN1uJbQ4mib0
Rxh89ExD788lM0WOfWBm7eS9VuYOtyeK0jl8nReYTlIYBvzIPYz8ml6tiyO5ocbJ1WOsw0Imdg0e
a0C8faTCbiOrkQ7STaFBAIEcq/FxL4GCWRmDzZHsChhtZ5WT72jNKz8YZbRr2wlLFdhFum37xuz6
m0SN0Uvn/0NsWEOdg4omezv05YF8bG0oubJFzZSaOzUkq+CD/ZhFjODH07tCiZ6uhwR2DtUhirpw
BlExZJQ4daMUD72du8FxpVoDlzb17ABVvczl9MKwCtMrg+NvWJZXEz0/+07qVagKgmj+/9X3Wwzc
SePEVkO4IfhoAbzpJf1IsE5SVo2gN79sHujKtBBvIEc+oaXbi7PyaJQGDjG7KGGDjCFxlXrUspcg
ETahlK4IIcF3g95l3xVHEjVkPxo75VQnjbpJKIUdukJSJbI6L4FGQK5NUg2Sak1wz8r+7a/mP4GS
TijGXHGg78mKeORzmEvnOKZmsIdfmcnf8g8J63fXwz7yY7nbhI6t2rhnpaPgkKAcqq2WEXCaNcLG
7FNMVdm/gmgmCKvC0q5UIJakStlVH386NMjMDyY4FKTWquafMa3z4Se1yByf7aLMz/I8hWbsPo9O
FjC3soM+2Is4m/Fxs3LbY8L+lH7snYDls+UHUqM8xbVR4kHEbdzSsRg0gohRAV3meGoGCuEaW+LF
el3QS2ztrSle9Qd7nGesd90+EKswfqQo1MQbnp7EZnVDI1YCsbgBKR5hUd1/ez9UifxDvabJJEWW
h/XqCFNkwFMWNuCq34LkTe9b+dhB2ghINQCp0k3yw6Kk0uEO4tfgQ+jfDU9NHvqtM0NeGl83LXEH
qP9/HyrWNHgkLbsNLeRWCVoB4DjnhIdu/obYkRAncrriYpC9RVCf9rilJ3bEhFDWrSiA+q8qKykz
ncbWcaLmv/i+Y+VWRBYhJrVQrcm2Z8+dLNcgGu2kw/V4wi3mwB/X7l4uZvaIPXIKqXgSS/KP6F8H
k+cAdUNrO7kZxGwHc81/4Pf7K5MgYEb+lYt3i5zgjvS6gWIbVX6Hk4nQ4aPGAhwfR5K0X7tsNRfU
RH2a3nKxNr8Gj8BaMV/Qk2e3QRh9MgPCMDmZ+VZEf2DZCEh09SNNS7ZagcB0sC76FeiTVjFbvNYt
DCsJ2OU+oa8+d5H+R3iROutIlfophUw9zstopkybuJy8WQ/qKQbjfrypQozspE3RIgPNrO9baj0g
Y8PZtnZdtHcebwywYOpjIYMqDseYJvYHF8X37s4CdT1BjpR/rrjK/QvnjwF35bZcEDmLMKRAlHEV
Enelz/4uQAcH583S5wYsBTFNC+IzUXvmhLG5okottXznVW0iRHioqqLgeFcsqvdIpI3rw5g7gGyV
Z7gHlUbjV8uneRXlGiiSWdryR4p5i2VG4vmQpR9HiX0/lampHGmjs8jE7j+isc/o3bR3zVdKLHqR
jk91wqLsy1uNeLeyZrI5IwsO8mSixydRSB/6wmkZ55L9ylHo+lEbOBXHq81HuSCjgkkZyOO3Fq0B
VoIexesAEb2zGY52epllxFOSDJLbMWhYKkPqJ1+YUK9gtaBc5aocu5YWpyX1D6IeylooYrsGMq8x
gdZiLzOQJS8z3Zzud2ZXNqp0DWYZdlJX3GvPMRy1Zd6Rf3ERTSfi4o0f4I8yq6WXefAB5LWvudM2
tGvhe5Bh2+rUfQZQwxBkVpYZ1FYi4onzbEV1o0PgEv10sorHzQTLM+ftNMeQnOGb1hg5YUiuxWhR
aUvj7Wvm1ZlP8kfKSn/zsLnfoslKD7sMmgb70ni2kDUQHI+sc0X0V7bAAx3fGEEpGiCfU45y3Y6n
qSswMi7trIu3gQhW1yXNFQeLFj0ViRyZc14pTSxfHpM2gmlXa/vecauyBFo5b8AiSBgEky6EelRb
qyFnKGQJL81Ugmy4wjebMBNx8HiurwG+LGd+TaQN7rIT61ckG60MeSL2f5e1PWpoA1tBn8AVjBZm
46SKJ/05QDi9AMMaYUeDIL3pxgC9ErsnOl+OnqWGCvWZPWUCiKCPrLQDIvVb1AxGbRKXDRMEYH7h
7zV0JE/Fc2C3JiPDuJRdMKjBj0cP4V+KkoNVt0i7jNvUBaj95QbISbMemVSnHs+QOtSmhgQST0fs
5U7n96dz260FM8vWrG5v4b1JHXqz4sGu6BbF7fRiJ9SkwKRlqEymy7m556j+F077s7cJojxUHYhd
nll4wqALbZjiV4CGJx95Sn15qjylsnxDuO4/n7Y3jjDgNwaa3pR1vzhhvAfM2CEOHgbx1lusyMA1
rLsDUNTDfuXwY7de1tvIRhfMoYdz87PTOoCUDmbVM+p3lPKDglePRAU6vblwDdDSVjcE/NGqxcv9
cUHxhuxRykyKtIfcxs9E+Vgb0dBn+NL6IClaiW7HepbLqAQxgSjO2Bs6qJ+2tFYhNKCl4HxXM8Go
Cuck/h5JdZXpnV28qx01MsVa/HefjT41TiK2uWhXsGEyAB6MHsNLVL6bNI2ie8+1qJoXJs321ZC9
Wr7A/8FcmdTjG+qcqtRK4ZfjQml7e8mEoKZQbxhzkQ8RZw38puXjj68WHMjiUc9O4qyfP0s7B9xb
LmhwUj2W7ITIwrzEaX5kllJy3B/7K0QtCer24CFz3kiXgENq+/OxYOCu2Z9LkTABJTuBvIun4NbH
qi+ksj/7tc8lyihHJGRdMvvwp4SWfrnfVro9HQ2VxuOwhmvOIMqqIS6bzMbly0W+aNB62Locaw1T
Sd8vlfWh6QkzYJ30NymCRHXuUOhf1FGhEOvXB5RtXuJnEHy2x3PqWNG6DlZNhEmsB/rGEKd3jN2H
W3GO7V9qId3l8SZknGbgiivns57Byq6C2wDctOW1qFPSSGntqRmmb36jdEyprBC8bxNDkSN1b6LW
iet19W7IrFrMEikd09rOkWz20JA8RRpEos+l0/Mt3DgD8X42QSZxbhXhbZQ2146sKUAvlip0GDS/
L7Roakd7w7J3jVc8V6KLarTfYsdjUTdzWXPRPl3HCQjnUfSnLjLq2igYxziqDQXnkM8FJP4ViYlk
Ttw3MQBE50i6PrEy4NzHPJUdNOjkjzHt24+OnPtsoo1nZmmmjfq7bcE9NNDSm4OWGrClm9jfrMmO
OCjf8VRV0U6DE84Er+Jl3c+SXHQbKPZ0/MG+h0H+56Hr7lIPCkmdJyOQcgkx+GOwbJYfAHWvjvMy
Gd8q+g0BnpPYDKyvpkS9naq0YBSvdc1l09EKvyo53/RoF7uzuC1O5pCkIbawWm4MkGVZ9fcxGsjo
jxxIskd3r45QoSZNFEqwaTNlEjY9ste0YJses5c5b6d4ASEyMmazh3Jys3yZOrK/GyLW9JtHnuZ2
7WrbX4KU/RTqZcjNGATdpviizlJuascF3bnmhmeuB0uqcgcrIn5/woEqhgPuJ/j2MWTovXHzejI1
0aHCwgK5HJTFykEDaXLuWILoTPEEeSHyfRUmK/glsHqrbD5p+KMrzgBG3missEPltN2vubfJXGeF
1g0vSfcCRFtTQ6jW/iZYOOM0aEAZfRmqwkJHsh71K0LkSEGMP/hmSGQ7yJfLDpg9jt8Wo7BLlUeP
nHMqe4CFpvt4p2A+N/oZUvwARPhWLAnpVm3eLhw4CSed/dQ+q0KnrGXXIktNaHKNwBPfHugtCH9Z
5dXRLEFTJfCAoR8rl0ucPoE1bG/ySxK3jpYMwgAQx0ONEiYk5gz4W0nL4dyL67bwgBPCXfwUsUOo
SXzqPeCF7c9mz0LH6Mpdl410I+Dlpdlet+C1VOpIaDwEjKFghcrKRd3e/wVRClnKdaSGVDYrZmAy
vDoOUvYsc6irkT81dqHf58tYrySB7jxa836YrAeCK9lm4uKuji0xA/abuSgcCK4A2FwXQ9n/aAnK
Gqf1CFAKqGse/oFGrz6ZmM+LWI2ql4tK1ZXuDcNus2xFqMmvgWzgSRCl2ay9vpNQdA9Pp5Xzp+px
TaJjiUfuEj6lflSrX2vIUry9dqR63YCKYOlt6xLncZArPB7BBsfYcragesO4Ky2KKB2VpGF230/e
MzclBM0uVnlSRItpP69g3a2K8v9i2QCjIOA/c3kBspHJcYdMM8tCjU0O53u1V9PRsOQ86hJs8rne
2jMZAk2WdZPNe5TkdL6Tt35+zPlhoXC2iC2nr1r80Ulo/AzoPDAehzt+uiczJyhYwHNrDCJosbvk
n59PUqJ7ZgCvrEefiE1c7IkHbsBEZ2NdGc58m92SD1DJgROY0kqfHhWIhXiywPEs9II74VyyjwgJ
iwLSZNv5NnZlwqDu5BxvJFVRixVfkweMdRtCiy5WDhmRvNg9IBqVjMZAPJecxkcPMmNrMtVQ2xXi
Ck5sUL7NIpnJf4POw8pa3jxscmPruC63AXvmq+CRDhFO6szUwPILaXVFGOr2gJbpFsJLcgWYtpRr
j8xg8aef5VMwOGiXmpSpgVMAXKyL+XZKSv97TXguNN1+ykrigvZZevBhZr754JTAGuj5Wo/zCmcK
Si4yAb3pqYI0lvdEJqqOxCE21VJy0Tr4YYPcL+r/TL/4epJ+Wpsj9U/rx0d5+KNvOb5flHCBp9si
O04w7cKf/7+ypSuZu1a4n+YLvi9x9/lQ9P1f5S0Mi5nCf9Iu32khqG2DDi0fY8N/CSFoRCH24ipK
dYy7TJJ9ozFic1AZ+5uG2gNl7rhl2FkO93JdF4PDV0vXKKjUziZIDnzTIriWD4xKrLjpVOEIRuhs
kYukxyeC6dDX8cMUd2NIkA8tKr95gM0kwCHDG1yf6YGGLFdrv+OKinytjOEeqmt1DZShlSTHx74/
KiaHEkSsvpcuzO/5SMS9MLBwegBCqWG9+6VTjSWcSojBM36Ss273UFjmZKu2r7q6vA9dCnxSu65d
UInfHBfgpf3DxIXJbF1bR+UpNsD7SSRvgN9Lj/t/VnDi8n9x67E8MGCmlgDXGpBZegYVadMrfufH
/zSiHV62xCbvv3haG7ZZqSO/gfBy29VEcYDNz4bhcxbFjZ2P8vAghYpIzYDci7wx3DRXonIBD52Z
BF0+o9RX2hgHv2Fr/phATZL2PLMAFKU6Hro3WBN14hgiBtnxDOEImuVou7NAto8E4c/7GbHwBbhb
YNvnLU3lIexeVbueRyCMetp4ytkxv04sXgX3VQYDZjusIvcxXZlcfnIz1s4Y+1GFUIhYVnH9wTwY
dq55wgxm8JDCL2+Qkc4ElPP1xSw5DicehrD363FuXEAHzgwOPECwuuwqBzBkIOucSc69rQBr7feM
ry2RuLqc/58MvqEyAndwNb7XDtwbNDkECeGp97VHg2gjNVAOaw43msAMmBlyQHlD4sfsnHqyePM+
XZuaistnp2Z/h44CMQooMk9PBNIHtjAlEymdiM9NVE7U8+YbjTtL8z/im168/DaTZ3LDHn1xxd/E
e9ly+npK8ihyFd004g7sJPdfs093wA/qkzQlDq6vWZQSAMZ3mSDAnq+5Ryy8l5KZeFc0m8Pajtvz
eVMtq5RViXTkf+k7iSqdFOs8FKb9Nbom7AX+dVoIdq5Wr/4Z7Ky7Afrh0piUZjzkG6OB6n/loI1Q
7HJuQ/DKl4E/bN+RUVI2U2sdVVU5mCKO2p4sy5sbqUT/NAyVzv0msLZu/X8l5yFY6oip81U4So57
unROlbets9UcHRruFx1txK316hiVWcDsMoBJKiepVPyUAHjHUKInFu8k1+vbd8sv1rUBJ7mnIxBK
RLStbY/ZL8NvbHJ+thSXY9mNw8bPCkyLvTHOJZbpiZdC0D60SgWhpCwb5qVEIRzKck8uCPDmoEYe
/JFgxIpnHKFjpX6e76YjTcBpbilOjhWyf6X8747mmC9wuXVFJBjdMS10UDhFMC+dwR03cpwHS2Pz
4uajTODmf/1wqu0aRpwN2P0D5wZtP0VLUlSupQjHVikXij4fCN9I7M7roVQ6vurgb+DzxZn2XvB8
Nk9Mty8RIy4+aRUhWFrUy75cnfs1PYN9Cdx5Y+CUtkB6Mi/BcYn3Nuqmq3MqlZVNbgiVzG1NZZ8a
Rmf4zTvV9DHwZglw7nNXdhDzp1NjKiudA9SP7+3610b8aceo57axmSrq6kugJDfiVuD6i+dPVp3m
OSxR3dmuhRK+NoYqzvejSB6jdEXZjgRBgWWESCGHrrzGvqxjWk6q+SCzxFPCPYzFjawrNhdlr657
5RknMHdclOGvQPkUy4xBlryZdcomcZA3MjzP/cG0VV/plljSG0Io9www3eNCVj+BellIPqkzEH6A
Yuxxqcm3XqvsH4wGX2XC/CYKLfte/sw3teuU7NWLMzZiVUMIF+johdKLrv2wvHqPAbGhPkYdkM2q
onKbFjnCcODN9jskc6kwZKImkp3y2KeGTFlrbtS2brhA62FP/SQlVdHhQDSVbDwd/I7ejIfmgMlC
pyEeLJtkNcvkVNg3dG2PZ/LNzyMJzW/U3hKbZKA4SBlRd8wqr4kxrQRFcTfoulJTREQTI/z7a89O
a1xbgd0vYgvS4wfKGLywvgDC25a1d3o5ves2phmsEaWxLiscuUCyFttD7NLFxqZEWPbKWsoAAkLT
zerJt01GVAFSAVurUajsJh0lxNk9ZpXuhEabS0ANVAos3HWAUg4TcTqlqrak9ysibM7tiV/2dtoa
fCD+CPITWlY5UMMJIbMONTrZlMZM87oqhg8auHGbWocAFJkMyNqu8Qh0oHzegNEB3P+1vAgEVH/Q
1e0JI6qMpXZyLHbHGTOz15uYLr4XKD+DezqC4C7+HnwlV8bgFzsx0n7U6QUgQpHsNLZ28xMaEyEZ
1X1odxSmKb5tSVNhTmMWrgaYtvH3DcdFPiGo0hkyFgizcCqbyWgPuoUvjb9VyFy6DUeGzFdg9/DD
Pq8GB+Ct/+Ug38JxH9HF7CW0KhPDaibqd3Akt52f1zov7L6chGL7YB0IlVbYDPtt8XABGD1erGu8
/4VCkL1iObIbmtD49uOEQJ7MSjQcDRU0JFSW4FzWgNIme27bbfn9T/p6namSRj9iKgJgSWYrSXXZ
h/CEkst0+LGH6LGgA9AA1iWB/+7TXuLVpD4ved0HKdswxxoOySeq3WZ9eizMK4Sb6ZDhz8b2X+/8
73DsiBvG3QLBBEyapKuEn6ICgqC8/YbEF8NEQv2dHeZzIRcMVHRnqRHnJ1QHVv+76ng/05iIeq1A
LEu+VawNOJPkZ0XgFeJOtYN7HLWjeCMKPvH2SBKz00lA1IHY6U5bgGjvCkk/hggo7OXSCCIoxNFS
j/eXTcqeP9eHopkQ6er3gRddxcuEBvvA4hrr6mTtdzclSLGotsLdjn+2biQQJKrgw4OUB70KTlD+
KxD4vHNwk7hWFZc9Csm79CUf5+l9ViTyJPotaQUM3V0DA0FCQI8O05Lu9Mes/G5xeU4LsNGkFWjk
YVtEFvrZN8ck88TBcotCuJ/Ixj+Gz3Bo/Z1gMFuLKmLm9oaF4w1WLq2Utlph8eBUTP0DzYPtaezr
/fqqXpwtW1iwhMZdIsu8+t3ShZ6VqKp4udnIBbWOls+/Uu6vsWsIdCa98rH5FValD+c/pvXvnoGS
k6wkn4FEJHghdRgaOVmk/+TSvvMQfmr2rerJrSN+EpegscldsuZI0azp7N0EqlBLp3z1ikMy4dKf
DOK+Z2+0Zbjb3JewNuX0gb1gp/+IlT0sS38brGJbcUYSTb9ud2AIT8uBv7ruwDh9R+wfTi6cro+x
GCICvdxyIdEUy4MwvW5FiuE0gr986oHEawukLQ/KktSAPNO9qdkd8TyAZIymN8zKBGDiUv+Mx8YX
swc7uvjd3WKtT04MaGq4LZj22lNYAwYtJOmJl3q43pe6LHrcyH40sjYp9rfJvF/pRHxteMBQ4LlF
16O4biCRZc6wO7/ScxIFyc2SvF6xwdOrJpx7ZMZYaCNDGiWTmkFoAPhdK+H/7S3h7Cs6hCJalyRk
7273WoA/j4PdaqXA3zJo395yd/1cwmuLJtQMaJZLHHleEqiJu3y8wTN0X6HmhIVIjVnPlqEyOQTo
l9/wfGTjTxtsPyV+oIGZSgbD8UkJzWmI3FY/q6W7gwuA7sh+4CEEHaVvm4PLsy102MrbyUg7IB8t
Jai4snfmeHcS3qp1+JBwkNkpi2nnnRV77UJU1/U/PJZK4oWLVPJcev03wlMO/9cTY32UPZgaBxZS
YUv1nczDpl6d7kMjMnDCbpMaY436f6br6JSdlBjKRgcX+Y8uYOnRFREFJm5gQGUtWrbWgxECCkN2
0tZXMOMfMdCw9qzG5X5x1gfoFpnAwIsZCyKVXEncmcZS3LiyMpqlQIGxBlCowcqaw6StPnOjnO0q
jVt3/vlmQNrCYqtP+EZvZa5HZM5eZ6wwo/LMi29LujH+9YO0QRE9APjk9R0AJwrtHyGyLWoROMqo
8orPk2jmM+zDeyeHewd+trExv4eHbxiu+W0lZutvVblyNz60k4TP7Qb1tGYoSb3VuH0gCgl1Nyik
s16tkq7K0nWYq0xZJ7e15hWKMY5YkdJlWHYxrtqf93is0E/zUhEFoqXrCD9i9RYrip81+KZqSwIr
hgiWIo7h5VJD7Z7zCLnOQuBXG51G3WpBUs+66TgIOzDe8D3oy+Ynd4WkK7GhriaZniPEwC4c9BV2
S/eX6BSLQvUXl9VvPwyKNhQadQAFI9hRTJ34e75YgENbC6g3Qqiy2WyoWp3p3QmhdwSejrCbcW6B
EK0LGcY8AuvWu3SXRz/O8oIHCrhHR0qE6vfv5Pw8Dx0xW/Cqglj1yd8hIc6aM/dSx1Mltd6pdgQU
MiZW9iNSufKkHMHEP7BmZhtQxnFAGsdwm/KbLqxes9nOr/lz9aMiZovygondYqzhGa1qBwaYZVe4
xQ/zcNq+qge8Gnw89BTOL8J2Z+X9UrobnAOIFGcT0/B1wC/4pDJ0F+YY0PaQptxCnS4yHNehYSlZ
TZohshysH1vLsZkjVgNfxaqGMQounC4UKkezoVD/LNSLzgnA41I/A7ZR6ncAzzACx4EdsqGL5ZDo
xLpAeal3pp3lJZg1tNPW6V203mv2VPAE8NXjnwMQYBJtYkgX6PAzHOnwpRU+6rkZM1VUiwsQk6Qw
44BvGsQjWuLLMumxARwDUgT/W2rwnHeUzhwcFlj3HFIUZQ18xPQj+VDQDDl8jmDqUfqQ+EP2vaxq
/f9MKeSXXrhSjKq1R370IlfhLZs2wyy5o7ZsgTH4pmeeuyk7siTNk9uBUs4p+lRm7tJktF0WTrRR
bQ70sIlNnOnZRY5c4qUYUbHgv+j34b0gboX/BhsxBbnyWg4jQA9eeCwsE8VcNxsrQPJCol1H2WlF
X5jnBqDp5z85WVHx9KqkxxMIhAmi/gLjknrbONPRMIXbdTa/b6CDj5c319Ht4Klxpk8QtP95SSvD
KzSORtTJwUPQBnN0ncL1GXI8ANPU4eIWSDhXetjkBeS+KJE3kd81vPrd/1xocD4I5WyCdRPsPi0G
NUTdpbkaDWu8Gq+pP65g+k0D3ocujG5JjXJiWhwwq94LCPe46w/BOppqr6ec+iyXCpwzjwq6xOTV
Xb9sFjlBb9HWH011HMihwi5M7Qq0JuC5AITfWwSX+qt6hEZhCfkv6oGgvoHae5bZ8CUWSvIOaWER
dOGKHqwrlZ77BdiPpD1bAQHnqcuiDGRHQElgy19wrQJ0z+zXH4msc4rmFFoV+fdOh0CK0tWhu4ef
t/6PjfGYay/v+hs8edOrjCX82Z4QaZ8uX/1OniNmHV6FTLs4Q8lUeoKjASFPmXA+xHE10CbsJkS/
U+GHSsc7c4+Av/STC4TY7Mf6eujujG/F0fiEqyUjAawiRYdnMyjE4bP+/jB3aMEj0c3PZhfpOkyF
D0bzIvJJzD/UbTlP/c6afjs2DtIXJjgv4beV22JKffCieAAZTqqiSIC9IFx5vv2FhSRydRJo1TV8
tm/2ijpvhnjDnQxBWV6bq8v0Ci0fkae46V5W1iP9hhux4CLgbfPfz5G1K5r/N1AvbntBuVjeb9yG
6ttwHCIU9xqB7ncKIpxfPIK0sD0bVQPXSzwMpntAmm13WWv4NAaGSn3P2O5j9AoZZ45XZwFn4uGi
jqKKp48b+g3Fu/Dy7u3sR6jwVTclwGKwfDQqjkJNi2m1hLmmtbKTuipcCB2G9eEYOcEfmY54+wRm
Hrscf6guxR4R6ZNb2YiMii2qa0Kw+7vkl0upVsnJPcgc+MvZthtv7ZhvEu4a8oF9LPL/txxc6crF
f2BgMGKMZ7eaIBMLKR6yu4deK70QiDSkAXUNvnKKL6hgIdTHsyIH4fxagudziWtwB7Vjj2Q8zL6h
a+qVyGeHxvyX1KH7wg+zOiPYJMHd5oQIYKgKADSG8Y+QLmYjRgcHP5gJUUMDTYOQ4N+5xmjZlk3q
ex4zL9+18AZ3knboS+9QEJGyqup9VvhGzqhY44yGMTpmIXkDOm93gmZKQsZUXv6jlIK81TdKLqRr
YhaOIVNey92g0tT3cv+ub/4LxRX6jd2CcI+7Xd7PWMYY2B689Bw6Tw92ra5D00NzXGER6zXfnMSM
1GIa7uTmoLK+U6Xd9Ur7es1hlctf9ARUEat4MqKnfx0rHIiZR2E6DL3sp3pG//xjLZ2pGXgEoDy4
RM0o3NoxH05DXbw0u0rolWMQCRZeJvrQpaDqpOY5SK5MrM/eJh/dUJee2M+f+fkgkfYIwqUM8CHt
YUp/9/50zZqCjcnmtHFRc1H37Mh1DmlGGhIRl9yUlg9mteQlbhhAcGuOjCAFuJbmPeOiDkL+8T9S
f6jlYydcUMv3aBIvf7M+SjPstXttx6AdKgK28JPer7SMJX6JSYbZW7FKBq/at8K/+UMBTixZsxYp
AIEoFrGdj6OaD4OFUgxEcpFoLV/KwOQD5qT9ln8q3uXQ+8cLJcwXEuzZ/a+GuPjZVSXaGCmrHlxd
Y5zr3gUTQf1j2jxuk6UFX4fEFrOu9kWMCm7Sr/0W3fSuFIxU9PVT5sCvJCOokc6//RFrhncZAubW
zP1YBZUf5fS5WZYH5ugvCa2UHr+Ld00DXxxu8eL1xnHsLxSQX1sgBl0mNLaOiXgRAM0zAtGBeVvf
/GrTxdl6H0AyFjimURhppvke+zoIdZx2/qErPWrsNSf9uqMG5CaPJNffE7WI7jCZDfp1tFxdUd/N
nEz4/0CUB7uf1JkOAAeXINhVU0rPQUVRuxk/qr38Yg0eW666r0gZUoYoUsmX4GSEdEToowbwQbK2
Wpux6j19xN6YgayJdy8byGRA58CFxkUPAPcIkWV8bp2T79YjeTnTvnuDkMHEfIoORPhI1UIiMwa5
bXLsQwMExS8QK/9+/BdtDMbl2LEpKNR7ByVyATEAv/EGEmeUlRs9NslUHC5n0Yp59jnhVQWiiP9u
zpUGJiOU01K7ty/bnCByPU9W0a6NqA2pK4UYUwajYNVjO4ZzSyZbdBJDnHkvH93079MWZwc8oiOv
4F4tiJhD2Kf/bfetptOYyElHITViqMdVhaOHJENr53NpyeUHfhDignof1lOxkMJ7/UgCwUYKcY+z
/tIJdoriSl3TN8YUGW/EaM0PhRTV/QtmKMm630QalkVDhc7fXBdOHgkNDNbx982rydVFBlJRGiMa
7WDkyNzUkFUwIEMf8r2xPPTQEUA3N+FrvsK5UA5bnyl+eK49t2E8HQRHN26lu5ftCLvsQ8SxMsse
ldGrasfWiC7LOd/OFNjEIKVr/VmCeewifkMJWInmw/PDfvTLnMdy0jLUsGbYNpVCHlKboAVYfJTx
D2MkKJnFgw00lKLlwrFab7st/9Vt/REbHdsmBx64lf5zpaHv60cVGnUkovhpP/m787vRhNS68Sxy
R+5sfgWwObGAIeIrH73yJWi91uM6Im1nrtGNLwbX0yA9L1c7IUBC82/LLFOrOaYdN215TyweaR7F
QTPlyK4ORI78+zrNhNQy4jQ8Y2rukn+xyuQm2fSwcDnQdeTyIxeQ9ZzLaeRoawD7DM1Udvc8SVgS
MFv+RSRZapQcPpT0iUmrcj7wuti2COixDMTwxZLQUqNOHTB3xopFGYMs5ZeD+2F+XMXIg9FGnyUf
NugY3mHj8QEIwwOdBRC2OAtKG6BuCKPE1N2jJMBAcVzZOD4c5l6w+HP4QnurMRbfE5iHYCRjCpFv
W/Q790GXLgpBX/FEgxLbjp/9aWIMO1SP79GvQi+tIwSk3a6pQoQaKZ152hi55Jydswh85rbhUZ4/
Ukd6dXgM8yM8FWZ5VCDc+d59S6B3FhqhgVYf+Oplqg0iWEVTY8khxatQDY9iPb1flwgS+dpPxIzn
nh1ujUNLQUh9KUawS95HsDF41bzzV1vLj4xJNyanRPWJKqQyKWawPUloLNAE5a/JtzWeuu0o4h6S
hfh94GCfTiQ6lZydgdLS5Sm2WEzhLFpgkQ91mujytX8159vvSJouPUZ/Oq6/sMefNpw+AKHiWcYD
7eklaRL1IzNq2906Zi+rTXA1vz8A18q86KfNT9QYoGx6mqvakaCQfmukHxUrZM25wMUoIPjFHWpB
wPOFbglQZLYZ9Sr0C0T/07EZdSS8/hXjg6d93444P/YhhdjaN5LrYoPI3yetfdXYRTqcTnHsx+5F
aqXGx1/f92KXdB4vZC3pJtUu5b931UeEl5nKtL4rxnGHO7zPTLfpYvBJ/4MND/cuLhDwqgRYs1YS
I9w53aMcbmuRErPM7bUNiSKyw+9LY0YJSgz/weE8klelNZd3ZYQTVO/ouKgPkEgQ3HHYUIyh6dOf
IrkirpyGI72sazRN9WWFEIqBge+CK+cOh7Ne7MZi9duKaSzfiWwWMcrdgelm8A6czsTpt+RVOzc+
ir/LF2ZZQx4D7QPdlEygluubpXjHkiPHwMGEQYVlKKrfd+C2TdKabXDl7tWzwhuVLsQY9U/QThsU
UQl03qfEj7gJ3gU9a7tqLFfbvHBADpJDemyhJE8iJ4j2M9+2N5YeV/RU2IJF/rd5w1/n1ro/SuS/
ZchKoUiW9Z/MTDXPuXJbjGvMYOh18WfQO2/C5eT8ZgEALbZAHABlzsWZ/NSgtBvTKYZPWO4lYUXl
4AZOJlhQ6Z2b/xbLQFV2yOPB6SORKUQwwy3DqTrOjxxohkJyCdGqbwkxYuWvKXX+/fWMcjd3TmUk
c/lIPc5vqu4Qj9ezJMWnR3ae/oqZdCc4HPyeEddMu9x/bbdfHwf+f+/zanq7kypDJx6JHljHp+fI
H9UqImZMUVGqkP2+3LA1a3DpM0xQgvEmcUnTYdXH3G6WolJcKkNxPI3G/NqAZPz5QYV7AvoOgQn1
scAq3yhjQXsk0pVeAds5++NZqFzZkQvbzXi+sE+pErbL/ZuOs5wgdKqvT2CsoZCabRY2GCVjPXRh
EAt0PSPpofHEVrbF5jj+UbuYUIm4jr35X4Wt03l70kCKILy5xMjCGgbtjup6i43ylCo2qlVpMLZ6
wf34gNKcZTkjCYeJ+WTU6AOzePW0j0+DoJ5KqzW3KGF7j2A9lu1ScZEYUAC+SGR8ZvG+JSiLepbj
vhPwcDGQA7ps7jOhgJ/zUP7qJzTekijsfZ/acGCPQDvU0y4IMzCyUQYBP3K7PHUZOxzanu0AkLWi
/wR0l8izadg3/RAAAJEEYqHVoYW5nZsSzkL647OuV98Q3Z+ZvLdzS53eKubRKi6saikPmWFIAeYP
sRZmRYAb1edHv9h8t2FH+bCjxt9/VTqgBQJ/8tc+8tbuLwvbKB/4B8UlrCbF2hTfOa+BfJVrfzXm
chzZVB2qmR3T4PyqkDzAAAOYy26ZIXcjMlRqJzl0b8dmc5z6aMQ3YUXr2hoON5qaCaQj5eb80eou
QSIToEtYrUxwIO4D3K33DZe9BqlZ6IYYTn3CFzcEGCWClv3Jub/q1PF1nJvfkoCWroSccMZiU6wM
4XSr/4WTvleCeevCNRHrcBrRj2cqizZ1kBnZ9p4zva5SL5s8nF5C1U9Gd8yWE2o2vMELxDYIhXgg
i2jMjE2fRyoCWxARNmXX4Pvy/WYJl8lFu20JKSaxV/45tR+gS83eqle49xlQE46XlaI+kc7JWgff
LUVE8hw6TQzi8epoZOh0uUJ8sDU62lrlfZINFLceQmuZU3ebLbt6riaJH3eq/HVgEWLV9j9xlGcm
2rq60fPIlTfCMKvQEr64Fwmnr5wOXEnZwT1dvLMAgasDFJ+bIs0dPgJR5jiCpvswd+ZTPsmLtg7o
IilYIpBWMO/lW8X1Upj1inslFci8NWCoJ7cT6jHLYLw+x0jdj6c6rh9efJ11V5Pypaf9iWan6rPd
ejVPS0oCXYxO7gaIhVp167r+vK/0QHUop4mjpn4nmIeeFws33r4vx1aHCbRcWwAIQNr3SUdmpWmF
09aWLEecm1z63u6CiUm7NWo/IziZ/TCkYlc3Aqk61Z+SE5CmjaKFrdxc6ZSJaxobwURs+k1Cw/C8
ZBusvTPoEDv7Y19cGzKfI4fLUlqsEnoGt6GOYZT1Z1bod4WkhhWyBWWU3Qeg6ZODn/xn170tI4QB
rycU8ebL3xExQfN4Qddv8PLeCKuDZdg2JE4lYhXycw/pKBDtD6IdUJrDRjMKhstBd+zibHX6VFWf
OPnSszJcIw1wvdfsjkxY/drRm+rZpOXNi0P/W8dv6bomwmoQGZwRtACfvc3vk6UGmL4n/sW0A0dW
lk5GIaKfKSBk1Q36gNfuDLItqRNcdotNf1sWwTuZv0n7hSJMiovNmdCII+brUN0pTOHK/Clt2q1A
wSpQniT71srHV5FYEazIL93b5ORbL3KJ6piyvJ/KZ7yLWMU8fquXL8T4UTAHe+Mr6uace8WAMlyX
ICUoqslDHoMmc8nz9qKjzO8GnQBkVFdRX/0nNPwlTG0U5MRsuKph3HQ/kyuPbKHTCkqEmTVXWJUi
pSZVV591eXyo4N5uvjcR51S+Yg4Mcik+XNyUb3OoDPKZ8pWJvX1tKrp9GIK8reQ6iItWU/viO0Xq
/zf9ZhXRIHKL6jAujJiE5vmVijo4i6R06pfLiIaITT/2+GAhH5xFGXnfdyDg9HxI/9IDI2SBd7oA
G/DQ1PshGJhNbHRFLfjp0tpxaFAU2uiqZK5DI8ypSNUhn20r972ZOAc8QzZuVz7gEi6ktk5wG3dS
qwsz30wyILcykaqJNz7wgWfn4h0uhAaLo8Y+QOCPvW1F5TwrYaqXVtOlvd8b9FM5D+H7CLLO19r4
+9Tdi666+b7jqm3Fb78VKso2RvUorqlfaqMYWVcD+VqcAtO8/ADjCNkd3CJNY+YGMcCPZaedu90B
6ZTtqCIhlcBNLAyvW54QmpMLmba7ZgobmoRf5lWRMTFT5zx3ItS/Zjt822i/TucvOmY/OdEb2qxn
69CQECTOW5x+s9Ya7vlk6pqN1HRaymuOF0EjdL/Qamb63W8dNsO0Q4i4kOs5U/uMRtXy8p7cl3+G
rxDg9HSFj5OtrN/GJ4dywYV8Z95DLFatYaz9lg0Klc6WPvjAMORICgPzKnWMxX3BLN6AiBmEc7I8
hE7hvaUKSBYcv0VJCXH9NcUBMNxXCOjqAnJmrV94aHv8uUaQj8c8ZHHzjtQo+FxJUSK7g6KHAZu3
9Ta7eZMu/Ooteje+XuGwmzu59xZXOU3ojyiUuDDg8XYpsBXWQM5bPfOatu98mxEyrAeq9bABRNjr
yFxPwxg2gQqG4yxhJ7WUwkL8E9SMoQHn/Iby0HLxVjJO1zWNMT7QFo3DnHwGFrQKqwfFC83iLj7h
KRzBcA9PAn/1/ljaJA5cK9h/it7cqtuwn5TVvzY6mOiKoLgkP8eSh+nPIpPTL+5HNp0PS+/aGEEo
rVSJzfo6E37AyEHVF+jt0JHEm2Ve1Vxl7mDzM9TwFdCgFHIESS+y02VI+Pg7aKW0ugTX9qzTBE5M
jt/jv7fiF86N104dgM64iGaMZEy0458dcw+BadDYRjyJxFT3tRJkB/IXqk2YzMaWR0/3aCrNNrHW
Jyz45E1C5bIluVoziOljveHERc3stF0FYA9re4C/mkpSpzOiMZjzZz36lAIk3Qdy1zlg5ct+nkOm
XtwJDS0dHd8qNXFZzZ6agf1KbjbyVSOQAoh6W9GoQ0pdR2vf6ZOBUgU499YO41feLvMTixbr3L8h
LdqCR8DC77oiYV1ol2M5qqQJn6yHym0ztbDKBSfoKB8ZlKD/tMoXZZ2LigeIYlR7VGI6Hw8LOHLJ
dL2oJ9uY8zEYKZn+X98vZUsYgJEuCQPvOWA66vFTX0hVpyFbwzxFEP6jwupuZG7RuntRIBtbTOIM
OuWAY7mdwBp5ZPvSArQxHHQK8pOfelVuvN/V4yeEaHAGHHYqqPy6NMwtB8nd1x9Pr+ePzp6o7Hv+
PWU6o5kEw6TuP0Q7GoH23P8tI0MADLmC/E2xBbFjkBb0dYZ+HJTepvvrqMlP5CFkfHw6J8bf2mCM
qM5tOWewtGKy9gjTWD8tj/NQ+/ZyaYjwKt/421SRR8k8m0obVtgPE0NGjW5vz2TW2aK/wPgimdG8
ujwRkoeKiqHC0CkjqtiichMx+LvSvuVVBmFGjFXxApvgeerd1pcDF2Nz0sD1H7HY2ds/TFVbr2aj
5Q3p3isGjU/hiGTbYe/lGdTJmnrPW1NCc17MDVioOFxHV+wG2iXeTnFpEXAsfGppB73uhwFV8E5E
RYw6fB+Olf4KcnXLNoOT24+Ir3uLJ0CSuy55K+eHJ5q6DflqE32zNaboSJS/rAoPcA5pV5T0pEU9
fJQrCPiA4Krx/utnr1a1Q8HGb59Qu5ETtfaLoZc1826Mx3i4u5wlY7Pgs5SYypnz4sSEynbB5LOB
g642AU8H9+rZU/0d94flkIuw5QrKV5F+ekLbOtr+0dNNDpwL2iCB4LUjeQ4mNFYk0RbYT86Xba+E
/BVnrHd8H+Xo5wRK1CcA7xo3sxKg3PIaIEn1/U4DDpwBlF4m6iuBZsHqhkR0duJ93kEu7UrxD4lQ
rPREcQCV5Xw+EOYDeK7A6jpkKM740WO1n7XAYTbLJnQOZWMJF8BcxRSHxuEOPV4QrDFo4/Yphhrn
ogzPZhw4kGPL2i58aWBAbvhceZzvL7MI0WZ9K8JXAelPayMJ4Q3FxO2kohZPj8y4Yp7s1LYuDDX8
EoM5FDI+r2Q2PuEGtc9V+zZmHvxZZIMlVcq53ucXZiuN2kvHBVSVFNwBDUk2SeCNYV6eJQdV0n32
QtLJodhIIM2w78VNGZ5tozw6UFZNsl+vs4dxIh3EBmObaL4PUvmwqvrsHDsXnWv/7qoQnm4lzNMt
PxWdoIL+lOPyyNMS3cDXbrLXqOYGfx+gnXJnDDTRgakRuDpeHAqIgjcc6eHlzJHo8CwUlGdYBlun
OGrkENp74NRszaaWP/5xLmMsMab0cj27p4PxUGqCW0JvgRlWJSYuBZep4HkRqjYvU//lNI4ZsX+m
yy7BE3QNohl5cGPSIpP+gLaK1cP8KSjsSi2JFUrYBmwC+DDUZ7K9acESOPsSlRm5nXwkF6StRCJE
AbHANmGcVjTIbnV5+3DHbFKQfhPX/0xfR9Jys4ykE9OvtBqJ7XNwMJecNtBBfMPP6HAxn7x/8+8T
wii4WqukhXBwYM7pimmDk2gthIeXLUyg1c/pLYzRyV32QHgh+uYFj+ychNmNaoNXGaNc5nXa8cxz
Ry86z7I3XJgGhTu1jz3GBe/UjMpv5kKzzJQGW1EBPmIzqFb8ZKcNRCGJnFuRU+JEO6OvDHViiFtv
8tDKKCYCpy4I1yI/2RYzMRuqJ+lOUC5B2P0WqcMAMaGTSZgMbgPecHD5yXg9ocl6Ex6VjrnwRNex
HKqNFsoGWwOV8scTFlIr5Tjf82ZiZzMsbHeQWF6/ujklxOQp67IUa/uAdIyyS+FJPrruF6bxB4oo
MtP/kItKVd+tiKmPj9+m9lB+v5GbTLGtUTtXvtaKomr1T4SrB4jcTRot2AFPo/uLWrp7zxnZiLVu
8++fa2gF87xCz6uYLk3TpLAWVLaOrN/CKXakx1NSZKJKUurb3VVQPGBCTF3WcaFOA+NKgW1gwT73
vzxAIatO4Kffyo6338StAibcGfS99dlPEAbyfQHkaiLzpQdKkTvISo7Z3IEpDpI3hrtbaXLEL23+
yl4Vdk73C1pBQhqGjT+W56+4M6chiV/LdAT9lxU094J0BirXCCQi5IHFn9oWus04rO8hlRDAEwpE
NyQZ/FYtN4MWzggS1rR+Zb89n57x5z16OMMVHTgMIzdkP4gprL1yMomZLZoPq5xK3Cwl78fY4GBi
tdhlCfyXI4BXioWjzXtUZx71JVzXxpmZSAeoqkObtX1eGpfND4qBjeD3uWgolULVJaRDSd+SDGJI
yBof90jSkAQP4X8Az7MieXvObn0HIjDJ5kVX/XhOj3uagJEjl6mMIU7wZ5+XUK5zniYVCjYY21q6
F235vSikGD6FT+wbA2M/vjbTD6FHEWbsAtPscJD9OGjk088JQsT4ExdF9V+lLDVazkQ+AAAKj/zE
qIpcvcnZ6nCV+bbx3F0ILL4Xh+A/Nd7bcj2Qqich4a/FA52YNLcMl9p04JmAKbLN0xig60ieeMeq
bn8Fz/+l+lk2AozYzh8YyiCLAtOgYw4Orn6I+VC6kG7wfRkaIVA8vNVr3oOw9I4o6z6YoffjvCDR
2zGwLelpavMjXL501rFIhaOSyR3DHKhyphl0/+aJ1o/86HJYHYEjJYPNphZIAjaxZAoMdhKCW/j7
RoYJUG5cz+yc8GfRIeNI+VtMTUQaDhnkuOylvYGvs/03glD08wQDHFtfJcLFnYgHNzL3nFet7kwe
LjBHPLBQfLq8fy9HebXgsNHBgEHuj8EXE/6foFkuYYeqK/P5B6gX2igd1K3Hz6eFumIp08i/nTJd
LtkDoWXd
`pragma protect end_protected

